// platform.v

// Generated using ACDS version 17.1 590

`timescale 1 ps / 1 ps
module platform (
		input  wire       button_0_external_connection_export, // button_0_external_connection.export
		input  wire       button_1_external_connection_export, // button_1_external_connection.export
		input  wire       button_2_external_connection_export, // button_2_external_connection.export
		input  wire       button_3_external_connection_export, // button_3_external_connection.export
		input  wire       button_4_external_connection_export, // button_4_external_connection.export
		input  wire       clk_clk,                             //                          clk.clk
		input  wire       reset_reset_n,                       //                        reset.reset_n
		output wire [6:0] sevseg0_external_connection_export,  //  sevseg0_external_connection.export
		output wire [6:0] sevseg_0_external_connection_export, // sevseg_0_external_connection.export
		output wire [6:0] sevseg_1_external_connection_export, // sevseg_1_external_connection.export
		output wire [6:0] sevseg_2_external_connection_export, // sevseg_2_external_connection.export
		output wire [6:0] sevseg_3_external_connection_export, // sevseg_3_external_connection.export
		output wire [6:0] sevseg_4_external_connection_export  // sevseg_4_external_connection.export
	);

	wire  [31:0] nios2_gen2_0_data_master_readdata;                          // mm_interconnect_0:nios2_gen2_0_data_master_readdata -> nios2_gen2_0:d_readdata
	wire         nios2_gen2_0_data_master_waitrequest;                       // mm_interconnect_0:nios2_gen2_0_data_master_waitrequest -> nios2_gen2_0:d_waitrequest
	wire         nios2_gen2_0_data_master_debugaccess;                       // nios2_gen2_0:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:nios2_gen2_0_data_master_debugaccess
	wire  [14:0] nios2_gen2_0_data_master_address;                           // nios2_gen2_0:d_address -> mm_interconnect_0:nios2_gen2_0_data_master_address
	wire   [3:0] nios2_gen2_0_data_master_byteenable;                        // nios2_gen2_0:d_byteenable -> mm_interconnect_0:nios2_gen2_0_data_master_byteenable
	wire         nios2_gen2_0_data_master_read;                              // nios2_gen2_0:d_read -> mm_interconnect_0:nios2_gen2_0_data_master_read
	wire         nios2_gen2_0_data_master_write;                             // nios2_gen2_0:d_write -> mm_interconnect_0:nios2_gen2_0_data_master_write
	wire  [31:0] nios2_gen2_0_data_master_writedata;                         // nios2_gen2_0:d_writedata -> mm_interconnect_0:nios2_gen2_0_data_master_writedata
	wire  [31:0] nios2_gen2_0_instruction_master_readdata;                   // mm_interconnect_0:nios2_gen2_0_instruction_master_readdata -> nios2_gen2_0:i_readdata
	wire         nios2_gen2_0_instruction_master_waitrequest;                // mm_interconnect_0:nios2_gen2_0_instruction_master_waitrequest -> nios2_gen2_0:i_waitrequest
	wire  [14:0] nios2_gen2_0_instruction_master_address;                    // nios2_gen2_0:i_address -> mm_interconnect_0:nios2_gen2_0_instruction_master_address
	wire         nios2_gen2_0_instruction_master_read;                       // nios2_gen2_0:i_read -> mm_interconnect_0:nios2_gen2_0_instruction_master_read
	wire  [31:0] mm_interconnect_0_nios2_gen2_0_debug_mem_slave_readdata;    // nios2_gen2_0:debug_mem_slave_readdata -> mm_interconnect_0:nios2_gen2_0_debug_mem_slave_readdata
	wire         mm_interconnect_0_nios2_gen2_0_debug_mem_slave_waitrequest; // nios2_gen2_0:debug_mem_slave_waitrequest -> mm_interconnect_0:nios2_gen2_0_debug_mem_slave_waitrequest
	wire         mm_interconnect_0_nios2_gen2_0_debug_mem_slave_debugaccess; // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_debugaccess -> nios2_gen2_0:debug_mem_slave_debugaccess
	wire   [8:0] mm_interconnect_0_nios2_gen2_0_debug_mem_slave_address;     // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_address -> nios2_gen2_0:debug_mem_slave_address
	wire         mm_interconnect_0_nios2_gen2_0_debug_mem_slave_read;        // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_read -> nios2_gen2_0:debug_mem_slave_read
	wire   [3:0] mm_interconnect_0_nios2_gen2_0_debug_mem_slave_byteenable;  // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_byteenable -> nios2_gen2_0:debug_mem_slave_byteenable
	wire         mm_interconnect_0_nios2_gen2_0_debug_mem_slave_write;       // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_write -> nios2_gen2_0:debug_mem_slave_write
	wire  [31:0] mm_interconnect_0_nios2_gen2_0_debug_mem_slave_writedata;   // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_writedata -> nios2_gen2_0:debug_mem_slave_writedata
	wire         mm_interconnect_0_ram_s1_chipselect;                        // mm_interconnect_0:ram_s1_chipselect -> ram:chipselect
	wire  [31:0] mm_interconnect_0_ram_s1_readdata;                          // ram:readdata -> mm_interconnect_0:ram_s1_readdata
	wire  [11:0] mm_interconnect_0_ram_s1_address;                           // mm_interconnect_0:ram_s1_address -> ram:address
	wire   [3:0] mm_interconnect_0_ram_s1_byteenable;                        // mm_interconnect_0:ram_s1_byteenable -> ram:byteenable
	wire         mm_interconnect_0_ram_s1_write;                             // mm_interconnect_0:ram_s1_write -> ram:write
	wire  [31:0] mm_interconnect_0_ram_s1_writedata;                         // mm_interconnect_0:ram_s1_writedata -> ram:writedata
	wire         mm_interconnect_0_ram_s1_clken;                             // mm_interconnect_0:ram_s1_clken -> ram:clken
	wire         mm_interconnect_0_timer_0_s1_chipselect;                    // mm_interconnect_0:timer_0_s1_chipselect -> timer_0:chipselect
	wire  [15:0] mm_interconnect_0_timer_0_s1_readdata;                      // timer_0:readdata -> mm_interconnect_0:timer_0_s1_readdata
	wire   [2:0] mm_interconnect_0_timer_0_s1_address;                       // mm_interconnect_0:timer_0_s1_address -> timer_0:address
	wire         mm_interconnect_0_timer_0_s1_write;                         // mm_interconnect_0:timer_0_s1_write -> timer_0:write_n
	wire  [15:0] mm_interconnect_0_timer_0_s1_writedata;                     // mm_interconnect_0:timer_0_s1_writedata -> timer_0:writedata
	wire         mm_interconnect_0_sevseg0_s1_chipselect;                    // mm_interconnect_0:sevSeg0_s1_chipselect -> sevSeg0:chipselect
	wire  [31:0] mm_interconnect_0_sevseg0_s1_readdata;                      // sevSeg0:readdata -> mm_interconnect_0:sevSeg0_s1_readdata
	wire   [1:0] mm_interconnect_0_sevseg0_s1_address;                       // mm_interconnect_0:sevSeg0_s1_address -> sevSeg0:address
	wire         mm_interconnect_0_sevseg0_s1_write;                         // mm_interconnect_0:sevSeg0_s1_write -> sevSeg0:write_n
	wire  [31:0] mm_interconnect_0_sevseg0_s1_writedata;                     // mm_interconnect_0:sevSeg0_s1_writedata -> sevSeg0:writedata
	wire         mm_interconnect_0_sevseg_0_s1_chipselect;                   // mm_interconnect_0:sevSeg_0_s1_chipselect -> sevSeg_0:chipselect
	wire  [31:0] mm_interconnect_0_sevseg_0_s1_readdata;                     // sevSeg_0:readdata -> mm_interconnect_0:sevSeg_0_s1_readdata
	wire   [1:0] mm_interconnect_0_sevseg_0_s1_address;                      // mm_interconnect_0:sevSeg_0_s1_address -> sevSeg_0:address
	wire         mm_interconnect_0_sevseg_0_s1_write;                        // mm_interconnect_0:sevSeg_0_s1_write -> sevSeg_0:write_n
	wire  [31:0] mm_interconnect_0_sevseg_0_s1_writedata;                    // mm_interconnect_0:sevSeg_0_s1_writedata -> sevSeg_0:writedata
	wire         mm_interconnect_0_sevseg_1_s1_chipselect;                   // mm_interconnect_0:sevSeg_1_s1_chipselect -> sevSeg_1:chipselect
	wire  [31:0] mm_interconnect_0_sevseg_1_s1_readdata;                     // sevSeg_1:readdata -> mm_interconnect_0:sevSeg_1_s1_readdata
	wire   [1:0] mm_interconnect_0_sevseg_1_s1_address;                      // mm_interconnect_0:sevSeg_1_s1_address -> sevSeg_1:address
	wire         mm_interconnect_0_sevseg_1_s1_write;                        // mm_interconnect_0:sevSeg_1_s1_write -> sevSeg_1:write_n
	wire  [31:0] mm_interconnect_0_sevseg_1_s1_writedata;                    // mm_interconnect_0:sevSeg_1_s1_writedata -> sevSeg_1:writedata
	wire         mm_interconnect_0_sevseg_2_s1_chipselect;                   // mm_interconnect_0:sevSeg_2_s1_chipselect -> sevSeg_2:chipselect
	wire  [31:0] mm_interconnect_0_sevseg_2_s1_readdata;                     // sevSeg_2:readdata -> mm_interconnect_0:sevSeg_2_s1_readdata
	wire   [1:0] mm_interconnect_0_sevseg_2_s1_address;                      // mm_interconnect_0:sevSeg_2_s1_address -> sevSeg_2:address
	wire         mm_interconnect_0_sevseg_2_s1_write;                        // mm_interconnect_0:sevSeg_2_s1_write -> sevSeg_2:write_n
	wire  [31:0] mm_interconnect_0_sevseg_2_s1_writedata;                    // mm_interconnect_0:sevSeg_2_s1_writedata -> sevSeg_2:writedata
	wire         mm_interconnect_0_sevseg_3_s1_chipselect;                   // mm_interconnect_0:sevSeg_3_s1_chipselect -> sevSeg_3:chipselect
	wire  [31:0] mm_interconnect_0_sevseg_3_s1_readdata;                     // sevSeg_3:readdata -> mm_interconnect_0:sevSeg_3_s1_readdata
	wire   [1:0] mm_interconnect_0_sevseg_3_s1_address;                      // mm_interconnect_0:sevSeg_3_s1_address -> sevSeg_3:address
	wire         mm_interconnect_0_sevseg_3_s1_write;                        // mm_interconnect_0:sevSeg_3_s1_write -> sevSeg_3:write_n
	wire  [31:0] mm_interconnect_0_sevseg_3_s1_writedata;                    // mm_interconnect_0:sevSeg_3_s1_writedata -> sevSeg_3:writedata
	wire         mm_interconnect_0_sevseg_4_s1_chipselect;                   // mm_interconnect_0:sevSeg_4_s1_chipselect -> sevSeg_4:chipselect
	wire  [31:0] mm_interconnect_0_sevseg_4_s1_readdata;                     // sevSeg_4:readdata -> mm_interconnect_0:sevSeg_4_s1_readdata
	wire   [1:0] mm_interconnect_0_sevseg_4_s1_address;                      // mm_interconnect_0:sevSeg_4_s1_address -> sevSeg_4:address
	wire         mm_interconnect_0_sevseg_4_s1_write;                        // mm_interconnect_0:sevSeg_4_s1_write -> sevSeg_4:write_n
	wire  [31:0] mm_interconnect_0_sevseg_4_s1_writedata;                    // mm_interconnect_0:sevSeg_4_s1_writedata -> sevSeg_4:writedata
	wire  [31:0] mm_interconnect_0_button_0_s1_readdata;                     // button_0:readdata -> mm_interconnect_0:button_0_s1_readdata
	wire   [1:0] mm_interconnect_0_button_0_s1_address;                      // mm_interconnect_0:button_0_s1_address -> button_0:address
	wire  [31:0] mm_interconnect_0_button_1_s1_readdata;                     // button_1:readdata -> mm_interconnect_0:button_1_s1_readdata
	wire   [1:0] mm_interconnect_0_button_1_s1_address;                      // mm_interconnect_0:button_1_s1_address -> button_1:address
	wire  [31:0] mm_interconnect_0_button_2_s1_readdata;                     // button_2:readdata -> mm_interconnect_0:button_2_s1_readdata
	wire   [1:0] mm_interconnect_0_button_2_s1_address;                      // mm_interconnect_0:button_2_s1_address -> button_2:address
	wire  [31:0] mm_interconnect_0_button_3_s1_readdata;                     // button_3:readdata -> mm_interconnect_0:button_3_s1_readdata
	wire   [1:0] mm_interconnect_0_button_3_s1_address;                      // mm_interconnect_0:button_3_s1_address -> button_3:address
	wire  [31:0] mm_interconnect_0_button_4_s1_readdata;                     // button_4:readdata -> mm_interconnect_0:button_4_s1_readdata
	wire   [1:0] mm_interconnect_0_button_4_s1_address;                      // mm_interconnect_0:button_4_s1_address -> button_4:address
	wire         mm_interconnect_0_rom_s1_chipselect;                        // mm_interconnect_0:rom_s1_chipselect -> rom:chipselect
	wire  [31:0] mm_interconnect_0_rom_s1_readdata;                          // rom:readdata -> mm_interconnect_0:rom_s1_readdata
	wire         mm_interconnect_0_rom_s1_debugaccess;                       // mm_interconnect_0:rom_s1_debugaccess -> rom:debugaccess
	wire   [9:0] mm_interconnect_0_rom_s1_address;                           // mm_interconnect_0:rom_s1_address -> rom:address
	wire   [3:0] mm_interconnect_0_rom_s1_byteenable;                        // mm_interconnect_0:rom_s1_byteenable -> rom:byteenable
	wire         mm_interconnect_0_rom_s1_write;                             // mm_interconnect_0:rom_s1_write -> rom:write
	wire  [31:0] mm_interconnect_0_rom_s1_writedata;                         // mm_interconnect_0:rom_s1_writedata -> rom:writedata
	wire         mm_interconnect_0_rom_s1_clken;                             // mm_interconnect_0:rom_s1_clken -> rom:clken
	wire         irq_mapper_receiver0_irq;                                   // timer_0:irq -> irq_mapper:receiver0_irq
	wire  [31:0] nios2_gen2_0_irq_irq;                                       // irq_mapper:sender_irq -> nios2_gen2_0:irq
	wire         rst_controller_reset_out_reset;                             // rst_controller:reset_out -> [button_0:reset_n, button_1:reset_n, button_2:reset_n, button_3:reset_n, button_4:reset_n, irq_mapper:reset, mm_interconnect_0:nios2_gen2_0_reset_reset_bridge_in_reset_reset, nios2_gen2_0:reset_n, ram:reset, rom:reset, rst_translator:in_reset, sevSeg0:reset_n, sevSeg_0:reset_n, sevSeg_1:reset_n, sevSeg_2:reset_n, sevSeg_3:reset_n, sevSeg_4:reset_n, timer_0:reset_n]
	wire         rst_controller_reset_out_reset_req;                         // rst_controller:reset_req -> [nios2_gen2_0:reset_req, ram:reset_req, rom:reset_req, rst_translator:reset_req_in]

	platform_button_0 button_0 (
		.clk      (clk_clk),                                //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),        //               reset.reset_n
		.address  (mm_interconnect_0_button_0_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_button_0_s1_readdata), //                    .readdata
		.in_port  (button_0_external_connection_export)     // external_connection.export
	);

	platform_button_0 button_1 (
		.clk      (clk_clk),                                //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),        //               reset.reset_n
		.address  (mm_interconnect_0_button_1_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_button_1_s1_readdata), //                    .readdata
		.in_port  (button_1_external_connection_export)     // external_connection.export
	);

	platform_button_0 button_2 (
		.clk      (clk_clk),                                //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),        //               reset.reset_n
		.address  (mm_interconnect_0_button_2_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_button_2_s1_readdata), //                    .readdata
		.in_port  (button_2_external_connection_export)     // external_connection.export
	);

	platform_button_0 button_3 (
		.clk      (clk_clk),                                //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),        //               reset.reset_n
		.address  (mm_interconnect_0_button_3_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_button_3_s1_readdata), //                    .readdata
		.in_port  (button_3_external_connection_export)     // external_connection.export
	);

	platform_button_0 button_4 (
		.clk      (clk_clk),                                //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),        //               reset.reset_n
		.address  (mm_interconnect_0_button_4_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_button_4_s1_readdata), //                    .readdata
		.in_port  (button_4_external_connection_export)     // external_connection.export
	);

	platform_nios2_gen2_0 nios2_gen2_0 (
		.clk                                 (clk_clk),                                                    //                       clk.clk
		.reset_n                             (~rst_controller_reset_out_reset),                            //                     reset.reset_n
		.reset_req                           (rst_controller_reset_out_reset_req),                         //                          .reset_req
		.d_address                           (nios2_gen2_0_data_master_address),                           //               data_master.address
		.d_byteenable                        (nios2_gen2_0_data_master_byteenable),                        //                          .byteenable
		.d_read                              (nios2_gen2_0_data_master_read),                              //                          .read
		.d_readdata                          (nios2_gen2_0_data_master_readdata),                          //                          .readdata
		.d_waitrequest                       (nios2_gen2_0_data_master_waitrequest),                       //                          .waitrequest
		.d_write                             (nios2_gen2_0_data_master_write),                             //                          .write
		.d_writedata                         (nios2_gen2_0_data_master_writedata),                         //                          .writedata
		.debug_mem_slave_debugaccess_to_roms (nios2_gen2_0_data_master_debugaccess),                       //                          .debugaccess
		.i_address                           (nios2_gen2_0_instruction_master_address),                    //        instruction_master.address
		.i_read                              (nios2_gen2_0_instruction_master_read),                       //                          .read
		.i_readdata                          (nios2_gen2_0_instruction_master_readdata),                   //                          .readdata
		.i_waitrequest                       (nios2_gen2_0_instruction_master_waitrequest),                //                          .waitrequest
		.irq                                 (nios2_gen2_0_irq_irq),                                       //                       irq.irq
		.debug_reset_request                 (),                                                           //       debug_reset_request.reset
		.debug_mem_slave_address             (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_address),     //           debug_mem_slave.address
		.debug_mem_slave_byteenable          (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_byteenable),  //                          .byteenable
		.debug_mem_slave_debugaccess         (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_debugaccess), //                          .debugaccess
		.debug_mem_slave_read                (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_read),        //                          .read
		.debug_mem_slave_readdata            (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_readdata),    //                          .readdata
		.debug_mem_slave_waitrequest         (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_waitrequest), //                          .waitrequest
		.debug_mem_slave_write               (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_write),       //                          .write
		.debug_mem_slave_writedata           (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_writedata),   //                          .writedata
		.dummy_ci_port                       ()                                                            // custom_instruction_master.readra
	);

	platform_ram ram (
		.clk        (clk_clk),                             //   clk1.clk
		.address    (mm_interconnect_0_ram_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_ram_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_ram_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_ram_s1_write),      //       .write
		.readdata   (mm_interconnect_0_ram_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_ram_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_ram_s1_byteenable), //       .byteenable
		.reset      (rst_controller_reset_out_reset),      // reset1.reset
		.reset_req  (rst_controller_reset_out_reset_req),  //       .reset_req
		.freeze     (1'b0)                                 // (terminated)
	);

	platform_rom rom (
		.clk         (clk_clk),                              //   clk1.clk
		.address     (mm_interconnect_0_rom_s1_address),     //     s1.address
		.debugaccess (mm_interconnect_0_rom_s1_debugaccess), //       .debugaccess
		.clken       (mm_interconnect_0_rom_s1_clken),       //       .clken
		.chipselect  (mm_interconnect_0_rom_s1_chipselect),  //       .chipselect
		.write       (mm_interconnect_0_rom_s1_write),       //       .write
		.readdata    (mm_interconnect_0_rom_s1_readdata),    //       .readdata
		.writedata   (mm_interconnect_0_rom_s1_writedata),   //       .writedata
		.byteenable  (mm_interconnect_0_rom_s1_byteenable),  //       .byteenable
		.reset       (rst_controller_reset_out_reset),       // reset1.reset
		.reset_req   (rst_controller_reset_out_reset_req),   //       .reset_req
		.freeze      (1'b0)                                  // (terminated)
	);

	platform_sevSeg0 sevseg0 (
		.clk        (clk_clk),                                 //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),         //               reset.reset_n
		.address    (mm_interconnect_0_sevseg0_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_sevseg0_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_sevseg0_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_sevseg0_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_sevseg0_s1_readdata),   //                    .readdata
		.out_port   (sevseg0_external_connection_export)       // external_connection.export
	);

	platform_sevSeg0 sevseg_0 (
		.clk        (clk_clk),                                  //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),          //               reset.reset_n
		.address    (mm_interconnect_0_sevseg_0_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_sevseg_0_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_sevseg_0_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_sevseg_0_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_sevseg_0_s1_readdata),   //                    .readdata
		.out_port   (sevseg_0_external_connection_export)       // external_connection.export
	);

	platform_sevSeg0 sevseg_1 (
		.clk        (clk_clk),                                  //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),          //               reset.reset_n
		.address    (mm_interconnect_0_sevseg_1_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_sevseg_1_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_sevseg_1_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_sevseg_1_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_sevseg_1_s1_readdata),   //                    .readdata
		.out_port   (sevseg_1_external_connection_export)       // external_connection.export
	);

	platform_sevSeg0 sevseg_2 (
		.clk        (clk_clk),                                  //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),          //               reset.reset_n
		.address    (mm_interconnect_0_sevseg_2_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_sevseg_2_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_sevseg_2_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_sevseg_2_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_sevseg_2_s1_readdata),   //                    .readdata
		.out_port   (sevseg_2_external_connection_export)       // external_connection.export
	);

	platform_sevSeg0 sevseg_3 (
		.clk        (clk_clk),                                  //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),          //               reset.reset_n
		.address    (mm_interconnect_0_sevseg_3_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_sevseg_3_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_sevseg_3_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_sevseg_3_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_sevseg_3_s1_readdata),   //                    .readdata
		.out_port   (sevseg_3_external_connection_export)       // external_connection.export
	);

	platform_sevSeg0 sevseg_4 (
		.clk        (clk_clk),                                  //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),          //               reset.reset_n
		.address    (mm_interconnect_0_sevseg_4_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_sevseg_4_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_sevseg_4_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_sevseg_4_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_sevseg_4_s1_readdata),   //                    .readdata
		.out_port   (sevseg_4_external_connection_export)       // external_connection.export
	);

	platform_timer_0 timer_0 (
		.clk        (clk_clk),                                 //   clk.clk
		.reset_n    (~rst_controller_reset_out_reset),         // reset.reset_n
		.address    (mm_interconnect_0_timer_0_s1_address),    //    s1.address
		.writedata  (mm_interconnect_0_timer_0_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_0_timer_0_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_0_timer_0_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_0_timer_0_s1_write),     //      .write_n
		.irq        (irq_mapper_receiver0_irq)                 //   irq.irq
	);

	platform_mm_interconnect_0 mm_interconnect_0 (
		.clk_0_clk_clk                                  (clk_clk),                                                    //                                clk_0_clk.clk
		.nios2_gen2_0_reset_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                             // nios2_gen2_0_reset_reset_bridge_in_reset.reset
		.nios2_gen2_0_data_master_address               (nios2_gen2_0_data_master_address),                           //                 nios2_gen2_0_data_master.address
		.nios2_gen2_0_data_master_waitrequest           (nios2_gen2_0_data_master_waitrequest),                       //                                         .waitrequest
		.nios2_gen2_0_data_master_byteenable            (nios2_gen2_0_data_master_byteenable),                        //                                         .byteenable
		.nios2_gen2_0_data_master_read                  (nios2_gen2_0_data_master_read),                              //                                         .read
		.nios2_gen2_0_data_master_readdata              (nios2_gen2_0_data_master_readdata),                          //                                         .readdata
		.nios2_gen2_0_data_master_write                 (nios2_gen2_0_data_master_write),                             //                                         .write
		.nios2_gen2_0_data_master_writedata             (nios2_gen2_0_data_master_writedata),                         //                                         .writedata
		.nios2_gen2_0_data_master_debugaccess           (nios2_gen2_0_data_master_debugaccess),                       //                                         .debugaccess
		.nios2_gen2_0_instruction_master_address        (nios2_gen2_0_instruction_master_address),                    //          nios2_gen2_0_instruction_master.address
		.nios2_gen2_0_instruction_master_waitrequest    (nios2_gen2_0_instruction_master_waitrequest),                //                                         .waitrequest
		.nios2_gen2_0_instruction_master_read           (nios2_gen2_0_instruction_master_read),                       //                                         .read
		.nios2_gen2_0_instruction_master_readdata       (nios2_gen2_0_instruction_master_readdata),                   //                                         .readdata
		.button_0_s1_address                            (mm_interconnect_0_button_0_s1_address),                      //                              button_0_s1.address
		.button_0_s1_readdata                           (mm_interconnect_0_button_0_s1_readdata),                     //                                         .readdata
		.button_1_s1_address                            (mm_interconnect_0_button_1_s1_address),                      //                              button_1_s1.address
		.button_1_s1_readdata                           (mm_interconnect_0_button_1_s1_readdata),                     //                                         .readdata
		.button_2_s1_address                            (mm_interconnect_0_button_2_s1_address),                      //                              button_2_s1.address
		.button_2_s1_readdata                           (mm_interconnect_0_button_2_s1_readdata),                     //                                         .readdata
		.button_3_s1_address                            (mm_interconnect_0_button_3_s1_address),                      //                              button_3_s1.address
		.button_3_s1_readdata                           (mm_interconnect_0_button_3_s1_readdata),                     //                                         .readdata
		.button_4_s1_address                            (mm_interconnect_0_button_4_s1_address),                      //                              button_4_s1.address
		.button_4_s1_readdata                           (mm_interconnect_0_button_4_s1_readdata),                     //                                         .readdata
		.nios2_gen2_0_debug_mem_slave_address           (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_address),     //             nios2_gen2_0_debug_mem_slave.address
		.nios2_gen2_0_debug_mem_slave_write             (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_write),       //                                         .write
		.nios2_gen2_0_debug_mem_slave_read              (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_read),        //                                         .read
		.nios2_gen2_0_debug_mem_slave_readdata          (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_readdata),    //                                         .readdata
		.nios2_gen2_0_debug_mem_slave_writedata         (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_writedata),   //                                         .writedata
		.nios2_gen2_0_debug_mem_slave_byteenable        (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_byteenable),  //                                         .byteenable
		.nios2_gen2_0_debug_mem_slave_waitrequest       (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_waitrequest), //                                         .waitrequest
		.nios2_gen2_0_debug_mem_slave_debugaccess       (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_debugaccess), //                                         .debugaccess
		.ram_s1_address                                 (mm_interconnect_0_ram_s1_address),                           //                                   ram_s1.address
		.ram_s1_write                                   (mm_interconnect_0_ram_s1_write),                             //                                         .write
		.ram_s1_readdata                                (mm_interconnect_0_ram_s1_readdata),                          //                                         .readdata
		.ram_s1_writedata                               (mm_interconnect_0_ram_s1_writedata),                         //                                         .writedata
		.ram_s1_byteenable                              (mm_interconnect_0_ram_s1_byteenable),                        //                                         .byteenable
		.ram_s1_chipselect                              (mm_interconnect_0_ram_s1_chipselect),                        //                                         .chipselect
		.ram_s1_clken                                   (mm_interconnect_0_ram_s1_clken),                             //                                         .clken
		.rom_s1_address                                 (mm_interconnect_0_rom_s1_address),                           //                                   rom_s1.address
		.rom_s1_write                                   (mm_interconnect_0_rom_s1_write),                             //                                         .write
		.rom_s1_readdata                                (mm_interconnect_0_rom_s1_readdata),                          //                                         .readdata
		.rom_s1_writedata                               (mm_interconnect_0_rom_s1_writedata),                         //                                         .writedata
		.rom_s1_byteenable                              (mm_interconnect_0_rom_s1_byteenable),                        //                                         .byteenable
		.rom_s1_chipselect                              (mm_interconnect_0_rom_s1_chipselect),                        //                                         .chipselect
		.rom_s1_clken                                   (mm_interconnect_0_rom_s1_clken),                             //                                         .clken
		.rom_s1_debugaccess                             (mm_interconnect_0_rom_s1_debugaccess),                       //                                         .debugaccess
		.sevSeg0_s1_address                             (mm_interconnect_0_sevseg0_s1_address),                       //                               sevSeg0_s1.address
		.sevSeg0_s1_write                               (mm_interconnect_0_sevseg0_s1_write),                         //                                         .write
		.sevSeg0_s1_readdata                            (mm_interconnect_0_sevseg0_s1_readdata),                      //                                         .readdata
		.sevSeg0_s1_writedata                           (mm_interconnect_0_sevseg0_s1_writedata),                     //                                         .writedata
		.sevSeg0_s1_chipselect                          (mm_interconnect_0_sevseg0_s1_chipselect),                    //                                         .chipselect
		.sevSeg_0_s1_address                            (mm_interconnect_0_sevseg_0_s1_address),                      //                              sevSeg_0_s1.address
		.sevSeg_0_s1_write                              (mm_interconnect_0_sevseg_0_s1_write),                        //                                         .write
		.sevSeg_0_s1_readdata                           (mm_interconnect_0_sevseg_0_s1_readdata),                     //                                         .readdata
		.sevSeg_0_s1_writedata                          (mm_interconnect_0_sevseg_0_s1_writedata),                    //                                         .writedata
		.sevSeg_0_s1_chipselect                         (mm_interconnect_0_sevseg_0_s1_chipselect),                   //                                         .chipselect
		.sevSeg_1_s1_address                            (mm_interconnect_0_sevseg_1_s1_address),                      //                              sevSeg_1_s1.address
		.sevSeg_1_s1_write                              (mm_interconnect_0_sevseg_1_s1_write),                        //                                         .write
		.sevSeg_1_s1_readdata                           (mm_interconnect_0_sevseg_1_s1_readdata),                     //                                         .readdata
		.sevSeg_1_s1_writedata                          (mm_interconnect_0_sevseg_1_s1_writedata),                    //                                         .writedata
		.sevSeg_1_s1_chipselect                         (mm_interconnect_0_sevseg_1_s1_chipselect),                   //                                         .chipselect
		.sevSeg_2_s1_address                            (mm_interconnect_0_sevseg_2_s1_address),                      //                              sevSeg_2_s1.address
		.sevSeg_2_s1_write                              (mm_interconnect_0_sevseg_2_s1_write),                        //                                         .write
		.sevSeg_2_s1_readdata                           (mm_interconnect_0_sevseg_2_s1_readdata),                     //                                         .readdata
		.sevSeg_2_s1_writedata                          (mm_interconnect_0_sevseg_2_s1_writedata),                    //                                         .writedata
		.sevSeg_2_s1_chipselect                         (mm_interconnect_0_sevseg_2_s1_chipselect),                   //                                         .chipselect
		.sevSeg_3_s1_address                            (mm_interconnect_0_sevseg_3_s1_address),                      //                              sevSeg_3_s1.address
		.sevSeg_3_s1_write                              (mm_interconnect_0_sevseg_3_s1_write),                        //                                         .write
		.sevSeg_3_s1_readdata                           (mm_interconnect_0_sevseg_3_s1_readdata),                     //                                         .readdata
		.sevSeg_3_s1_writedata                          (mm_interconnect_0_sevseg_3_s1_writedata),                    //                                         .writedata
		.sevSeg_3_s1_chipselect                         (mm_interconnect_0_sevseg_3_s1_chipselect),                   //                                         .chipselect
		.sevSeg_4_s1_address                            (mm_interconnect_0_sevseg_4_s1_address),                      //                              sevSeg_4_s1.address
		.sevSeg_4_s1_write                              (mm_interconnect_0_sevseg_4_s1_write),                        //                                         .write
		.sevSeg_4_s1_readdata                           (mm_interconnect_0_sevseg_4_s1_readdata),                     //                                         .readdata
		.sevSeg_4_s1_writedata                          (mm_interconnect_0_sevseg_4_s1_writedata),                    //                                         .writedata
		.sevSeg_4_s1_chipselect                         (mm_interconnect_0_sevseg_4_s1_chipselect),                   //                                         .chipselect
		.timer_0_s1_address                             (mm_interconnect_0_timer_0_s1_address),                       //                               timer_0_s1.address
		.timer_0_s1_write                               (mm_interconnect_0_timer_0_s1_write),                         //                                         .write
		.timer_0_s1_readdata                            (mm_interconnect_0_timer_0_s1_readdata),                      //                                         .readdata
		.timer_0_s1_writedata                           (mm_interconnect_0_timer_0_s1_writedata),                     //                                         .writedata
		.timer_0_s1_chipselect                          (mm_interconnect_0_timer_0_s1_chipselect)                     //                                         .chipselect
	);

	platform_irq_mapper irq_mapper (
		.clk           (clk_clk),                        //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),       // receiver0.irq
		.sender_irq    (nios2_gen2_0_irq_irq)            //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.clk            (clk_clk),                            //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
